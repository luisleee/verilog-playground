module d_ff (
    input wire clk,
    input wire rst_n,
    input wire d,
    output reg q
);

always @(posedge clk) begin
    if (!rst_n) begin
        q <= 1'b0;
    end else begin
        q <= d;
    end
end

endmodule
